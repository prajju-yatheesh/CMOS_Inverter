* Testbench for CMOS Inverter
.include cmos_inverter.spice

Vdd vdd 0 1.8
Vin in 0 PULSE(0 1.8 0 50p 50p 1n 2n)
Cl out 0 10f

X1 in out vdd 0 cmos_inv

.tran 0.1n 10n
.measure tran tPLH TRIG v(in) VAL=0.9 RISE=1 TARG v(out) VAL=0.9 RISE=1
.measure tran tPHL TRIG v(in) VAL=0.9 FALL=1 TARG v(out) VAL=0.9 FALL=1
.measure tran power AVG P(Vdd) FROM=0 TO=10n
.control
run
plot v(in) v(out)
.endc
.end
