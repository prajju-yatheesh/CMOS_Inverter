magic
tech sky130A
timestamp 1694352000
<< pmos >>
rect 0 0 2 1
<< nmos >>
rect 0 -2 2 -1
<< poly >>
rect 1 -2 1 1
<< metal1 >>
rect -1 -3 3 2
